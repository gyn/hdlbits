//
//
// https://hdlbits.01xz.net/wiki/Step_one
//
//

`default_nettype none

module top_module (
    output  one
);

    assign one = 1'b1;

endmodule