//
//
// https://hdlbits.01xz.net/wiki/Zero
//
//

`default_nettype none

module top_module (
    output  zero
);

    assign zero = 1'b0;

endmodule